library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity F2_1 is
    port 
    (
            
    );
end entity F2_1;

architecture rtl of F2_1 is
    
begin
    
    
    
end architecture rtl;