
module unsaved (
	clk_clk,
	reset_reset_n,
	entree_anemo_vitesse_vent);	

	input		clk_clk;
	input		reset_reset_n;
	input		entree_anemo_vitesse_vent;
endmodule
