  --Example instantiation for system 'Sopc_barre_2'
  Sopc_barre_2_inst : Sopc_barre_2
    port map(
      clk_adc_from_the_AvalonVerin_0 => clk_adc_from_the_AvalonVerin_0,
      cs_n_from_the_AvalonVerin_0 => cs_n_from_the_AvalonVerin_0,
      ledBabord_from_the_Gestion_boutons_0 => ledBabord_from_the_Gestion_boutons_0,
      ledSTBY_from_the_Gestion_boutons_0 => ledSTBY_from_the_Gestion_boutons_0,
      ledTribord_from_the_Gestion_boutons_0 => ledTribord_from_the_Gestion_boutons_0,
      out_bip_from_the_Gestion_boutons_0 => out_bip_from_the_Gestion_boutons_0,
      out_port_from_the_Leds => out_port_from_the_Leds,
      out_pwm_from_the_AvalonVerin_0 => out_pwm_from_the_AvalonVerin_0,
      out_pwm_from_the_Pwm_avalon_0 => out_pwm_from_the_Pwm_avalon_0,
      out_sens_from_the_AvalonVerin_0 => out_sens_from_the_AvalonVerin_0,
      BP_Babord_to_the_Gestion_boutons_0 => BP_Babord_to_the_Gestion_boutons_0,
      BP_STBY_to_the_Gestion_boutons_0 => BP_STBY_to_the_Gestion_boutons_0,
      BP_Tribord_to_the_Gestion_boutons_0 => BP_Tribord_to_the_Gestion_boutons_0,
      clk_0 => clk_0,
      data_in_to_the_AvalonVerin_0 => data_in_to_the_AvalonVerin_0,
      in_freq_anemometre_to_the_AvalonAnemo_0 => in_freq_anemometre_to_the_AvalonAnemo_0,
      in_port_to_the_Bouton => in_port_to_the_Bouton,
      reset_n => reset_n
    );


