  --Example instantiation for system 'mon_sopc_pwm'
  mon_sopc_pwm_inst : mon_sopc_pwm
    port map(
      out_port_from_the_Outputs => out_port_from_the_Outputs,
      out_pwm_from_the_Avalon_pwm_0 => out_pwm_from_the_Avalon_pwm_0,
      clk_0 => clk_0,
      in_port_to_the_Inputs => in_port_to_the_Inputs,
      reset_n => reset_n
    );


