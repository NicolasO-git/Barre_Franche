  --Example instantiation for system 'unnamed'
  unnamed_inst : unnamed
    port map(
      out_port_from_the_Leds => out_port_from_the_Leds,
      out_pwm_from_the_Pwm_avalon_0 => out_pwm_from_the_Pwm_avalon_0,
      clk_0 => clk_0,
      in_freq_anemometre_to_the_AvalonAnemo_0 => in_freq_anemometre_to_the_AvalonAnemo_0,
      in_port_to_the_Boutons => in_port_to_the_Boutons,
      reset_n => reset_n
    );


